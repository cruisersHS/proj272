// This is a simple test bench for the permutation block
//
`timescale 1ns/10ps

`include "tb_intf.sv"
`include "ps.sv"


module top();
reg clk,reset;
reg firstoutH;
reg [63:0] din;
reg [5:0] dix;	// data index for 1600 bits
reg errpos=0;

wire pushout;
reg stopout;
reg pushoutH;
wire [63:0] dout;
reg [63:0] doutH;
NOCI bif(clk,reset);


`protected
C-#0c:^eG@L_=1C^_T,/[IBe:F8^U&#.AR@22HYQ>^._S597#e11))C;2@/?dFPY
=IT=F@B]Q/eUZ&W)g6gGb7V8O)UDZZ(V<CGbP=PVT)8)=+9gdZN[7I&aQ3/HVU3.
KFY^2;.C=T2MV3G.U)F7DM3>_5[DbP,K__;[;RdD#;_FEa8>P^3;QK=01:c9R1C#
+D6Q6Tc24eD7@&QMOYL,@Td,e-QIZ&O=R,S]2Hc<JaJB:O?U._WELVISX\dFeK?1
aZ(-=5Y3=H.?f,93H60,JG8=/(G>F2NF+CZaLV0d=SQUEda^786P6IIF=gK?LO#_
1QK<RT2@RSGIY]0(3]Yg]H3/U^LZgQMTZbT1E=V.2(04IU49MXS,M>&0)RUfB-4D
5XK?PdW2?,;O>TIH6&T(fJV6bAJ&Y^]&4+=[4:6S206CWG9<c/KP9(e4/R)\)RAF
]H>:Nb0>.K9.,KW,c&\G4&a\4[5+0\ZRN8.6dG&4H?<Y4;J;C7KD3/6I/d,-5f>/
&09LYcV[YQX9;F8N,Q)@fMM>VgX>b9L?O7GI7(b21<GQI:=(KZgFRC1MBEg69>+<
9X\&7M(Z>;62S<W=I9&QBU9a]0Vd3^2E/=GK@-/S+)PA@]-T^ODHGeE\]>gSDNLC
)Z[,JJL6LdAF7BT([1)NAEP;E?5#I4(_X0\JJ7]5gP[;\cWcV7_NF=(RX\BFR)?V
68Zd-7_B^UJ+X0ALdF4^SBA4O9.XRKdXf)0B3)O0^NNI28QH[U&[3QA7@(VX5>O-
HEdTC[H2&1SdQQc5/4D76W8)IBcO<6K(gDQ3OWQ,6@)d@a?MTNS<[H;,S^,XaFf1
0D\EfJ>IRLMQeUH8ef,5E^RJYFIW>#UNT9K)\QG+<G7GN-Q?FeWBE[.QBB)c\aZ,
0X1=b\N;Og(#e6?]SOZ4;,25NI[#.\215f4-#FMEXHQV>X-Z><b;8;.7:\eaa9CM
CSUD_Q>8UZTE8T&VJ5B7,VL-eT[#M>L(9AD_B]2J[YE919d1JY<bXQ&/?KBgG\15
2SK&B6H\DU89LCBDWVPHTC5:(__DEefN>SL4=5P8NegDFeJ9ET/)#6MbHA4?^=R)
@2?BLX-aAJ)?4];gVgKMVc&g&_6I=X91TDCLJ[_]8=bJRXfBI:8bKW2HG[T5/M(J
_RbEM&R3X2H9X]#JaB:EOa=,H[6+J6UY(<(g=26CXC1/aVYHZ?&+Q\7;a@g]6caA
L+g7QcA<X=)Sa71,&MBZCQ8:g-=6<Z<)1,:C7F/A9aCJ5G:90],Yf@#FR:54Z\e]
O(5>baf<A.:_DbM(FYGdL4](=;#8:.?CXK:X?+]3+1Ub-[VZY)@]1W<&FY#L.Dd_
=3>0)S0+AOT5\B<PTL[IE^R.fS(DI_?\DUR]R+6.F998Q48UF#.gY@67(MGUDT98
,G3;&V=V21J[M3#B+:0E0N/=RNXSU&F4[a0.DTS/Q54#<P<]^O<]?_3OV3L@W]+H
.?O@?;G4M5SD=Y#S)4@\PX0>&7dDL)C].[J/N=HG^S,L.Ne6VK>_3/9]ZKdSS#g/
T5d)=K9eP#C(YM\\9bc)[a/M5HQ<?COTg]@E;D6@._X=Vf3d[5ITP?Eb&1A/XP,K
;3d]cVeBBO#6FJ?GJ,]R_L8?<CG)c-M^P]bS;/;?JaM2Lg(.f+aF-)gO)])FQB,Z
(8/_?>S.09;6d@=BEgWaIJ?F_Z_Y,/G_30:ON]7V-\8#2c=J:]Jb^ZE;N8N2A3dU
6#Yd5V)]aQ6#ZLaf4MV4T:67M/S-X;L)Y]PF#T@C6[?g?5]\[O@1EL)/g(8T638G
QS;]XMfALPQ;I;L>9V3N0=Z9BV:TfdEe^[(Yb5NeTRg;(&L4d<,KF?]_\=bBF#]2
1f@R@9B#dZ0@(-YB+Zc]D=8_#4_GBC,V).AF]77:#.B;S>,e/4X]7<9dC8)8#TEg
285eeQ89]:UATU4gB/AVNLTVdI8>XS3(;Q+WUd(L:B84(HI&;O0&<5P5#fb[dAOO
<+VSE//b^QMO:+R9W[aXeN<e,E\MFIOF_^a[2f&a>CHUI6Ad^gSaC#AWL?\PI//A
QB](?=9/)\/,_91Y;@(6-9Ig5,R.cD@b9BVET)-/dA[8V^P?\VJ\9:U>JH^bSD(N
,F6d_XW#C\<_8CEOYCC-]<8JG#b-TN]H64+YP?62HCA>C_aHLOMCEeOF,,G;^O5^
T];X2?bY537[bdBa=N4@HRCZ]NLAHSM/E+63,7URJOK^R(LOR4?EQ[#4\K/Ag?4)
eJF=CDTYH3M29K678--4#8(NSST^MNG=?:/,Va2^C-E]7A_C0^4Q[f1[A4#:I>L3
GP9U^U\U6fYF<RO^IZ^/#.Z1=)Q3OdLXV^F;4O?>+-APbHX)b<_g(HYG9&C?Db1f
QLX70b]D<a;aMfd]>,9g1700TLdf_2DLJ8)>/gaL<a^;8YJ1V.[LV>W5#K4,JNZ5
2/&WV9T=>_(JIfGeUKCgJW5/(7g8:J;P(J-+,P0Z,?;C0).BQaC]-@>dQOK2MRd)
7/2,E3LcH2X6T3@\^N:CVFJ=&._]S>6?eH2^&.?_,V3W?=db8&16;G..Y]?SS1JS
1g9bQL?\?BG<<:#1N4&[8^BYI?@OEE[<\a0dM&W,2IRWQ^HeMY<PHC4O;/1E?D-A
9LeVW8LG&;IJ^4IQQO/M/)KR0^&41e2^L>dI97U-/6>/SR7M^fN49UNTG5KC_B.d
Y>d03L5BD==&([&?<fAY3;MNeO5e]K3I5G_;;&+,G,3@@aaKR-^^?\;,[A]U;K.;
IgU)F@^eNZZ)SIP:#;@K(f)#LK.=ED#STT,\\/W8APZ4U\<499LO&58[V89AWPHf
,,;H,91,V02UfL.UR0-]6PXM_QLdI]JFXQc0O]-G1c)&B7T=Z#OJF<HI<]/gcEBB
NOR/CPDd\H=NIXFCb+DZE7.(IE:gDN48G=5a99/P+9I_\23TB+?F9c)7T03N=QbR
ZD:J?DKdZEF,A#X)XK=1=I]e:\d:]e:D\RC/;<Db@Rg7.L<C6Je\SFMcBeWI76+A
XG>-[Pg>5g:CVBB&(,,8+^2X[f<e5LWbR27H7=V-AI+/XaM#_/E1[5M2<325<<K+
QI@4.1:+K2H9A](8be3QI(F^/(AD.MdWE,Q&_bY1KK\gBI/9RO9+VC#=)<6LDFB4
9Z9HN9+<+?baTM(1I5>/(,Ne(K\2LMHV?<7LMM1?,I2MGSQJ@UL2Gc?e\,/2TD.6
0K@+c8DKa\,:#-a(XTX]HXcL<N/,4&<H[eJ4J^\9e6:[@?85Vd(KVE,Z/2G.bRd4
Og2d8)CJARHda.D93643.f4;J=VX6MN9NP[W#LY9NbAcSD7W.F6KU,]C(;f/1gBF
<J0b<,J.B1,5,X=523H08Le_Rcb1Fad?N@/L5E;a(.\O]>JbRKO><Vc5@..VZVKG
,N@[26DePM3W9>0^_9D]H7dB--I>M9DagMY2+]d&Q9a1a99@T2=O>_>._c&:.G;2
YZC\1+OHNgag,+-gF^@VX07N>>2:7;=42(Nf01f3QB4CQ]MVCZ_.1;JX]Lg.Kg=&
KG&9V0IA1+^@3#(F]-.PUNN6dEN1KLfUgIU6=CE0(QGf=,6b/;c2EB(PP]PXDFIT
]g1VR5#?[E&/RCQ:70>QV<--B)#HG1b34F_?WV8DT[Ca8c2].g:H_,;WQ[W6Q[P8
_)U[-7.Ica&@bfOH?fK)@Ga?\]HJ1_(^HDED/6F_R#+P#UQN2RB,B/bI<+:G:0W)
07+AY;@[EHg^GG_JXI#f/.(NGebb@^:7_;J4]JR?(9aScH\c)LM225;CH/:fZ;g.
P.,<=HE<XQaV\QTb;=8F^6Oc2cDZaL=BD#L.(#VD6N;9)218P?(S=4\+OP^a=@L+
2;.=/M#&Y(UM+2BPaV?:P(=YdSF32W5_P_6_SU[RZTcLOCbYUcM4Z;OELACBY&_-
;KOd9._aJ-eb@).GbdM;6^Q_&R2Z(XSG;PcH5==IBM;/H:=U><#;1b8gb&M?B+(9
X-F75>7OBb#MLOg8cB4,6F[:0dE0fCP&GY@XcQ#1PJ<NaPg2&<R4H+[5Z.;[]EW\
B[e/dZ)6X0/+I)]=+7V;:0bWSd:]Z.XI&<CR,B.M0,f<F3,YAM@bLGXA00M4[8PF
&:VB3_EDgL>T;fIF;Wa>GD(6ce+U??O@dJeZDa]VIFYZ7])&-J5aFFG;f+@S=a^a
fDccB7dEZO5.UEI(Oe,3YT@F,]?GUF=g?)8K+e;7T/P+67C<1K?dN,+-XVcA@2]5
a5Y\WKG<K4/)A/QJ2&E^)E^E/4[)TV6,?+F:5<(aKWSd@E:W-aa^]:KW1.;4?S9Z
6Le-d@D:373\^Ha(,fR,5-+KQ]V91;+HMJZ>\F+D1L@dW11M?H?2d;#/L+E4[D<,
Q?8eHY4XYMG@0)L/bB^PM[E01@8Ga&-fFOOdD3@@D_GZZ@Gc/g4^U_]1[3+[eU+1
&g@5Re6#>+T,HDRa,/Yd(PSF0<f&-Q?&XN._+2):CXYJ]Z_::Ve:ROHH,KdFJS5a
L?8YSWU2c_E7ECSQ4]\H<B#5g1e]Q/dQ6-45OeFR/IR1N5:@RCeQKdf,ON40M3HQ
0F2CTHQQI(2aW-ZK@geUZ#Me&8)E9GAA>T8PA\5<K:B^fX\UH@3LS;a>a]K2>g_&
AX>Y@g-?U(6a[6JPG1JC4AFE54X[0f][XV/C0?^Ke:c8C&CBLY=_8Kfc0d(=H&;N
L.K:HQ/QE,_;OQ_aJ]==g.QRFYFOZ+&I;#+Z[7Z:^)+\ILYMa_;>#:RZ1HJ2@bM/
6dTH0f_R]U+dc28(cN6@I=5M;I0e:<[:,CRS[D.E;;(H;2Y,STUV[.)6g8b(G9eE
./D&RUE=3Ca7aM_?IR#7]GF2,C3(++R9(2@&>TUS3]^3SIL)95K/7[3LN6I?QB&H
SA_@^@9LcI>\_?49dMR;g0SOW6K\#QETQUW?3=Uc/=d0UX^[=<L]_.M<[K@=I+g[
[POfB]K3]FG@/_952_?NbT(Q:AEg+GgPYA=3N6OSZcc9]@#4+^.2YG;]L)8e_OWg
OJK6,d9K@[Zb-5V@QZ30]UW?D@Z/\gP9JRf]R&F&a5-(>cFWWeVN>XJEf_GZ-^e(
@TJ.A?&QVb2g>Cfd+&[WGeT@6GG>R@)g]D+Qg,0:U]e92:99Z?U<]9c@A2S7CDAW
NOP?-Q?\H59WG90,FG[,SWX+@)<].)&/EEO;]2c/=X.]DKA6?@QgU-RWD&+EHU=]
g5[F3c#<#L25J7INQ#_2a+&/8]CBU>&MS][dB=>K@J==IGZ,7_e79bUP_)?2D1CG
Y>M\cZa#^RA,3UOA7gB=+a8_G12Y5/#X;Jc53-_;9ZS.)CXB,96:GFB.U=X9bgMQ
-^XI2/([.Pc>5\=LBPLgMR:,BL-QW)#NCA#b0?\gYV/4.eC@^Y@&@E/[.H9=/[#0
=+M\?EH([_-LCN<&S@ERbSQT1#18=:R;AO?aT5;,9]dc@9=>@(DfN/f-cRZ-UG;X
UAdVS.-/g,7V34+?BUd/K](628<]7.3eF+T@3\2HV-]GOME04B2UHG\H(3B:NbI,
FfbNB>4be_-)(#D@71(6FdD0J6;(:aXN(C_:Z+GecQ/^f?Y&7]BgP@6:eXJ+8N]W
93KH=KP;A;U.\f1(Rgf7WO#bM=c.(E]a_0/gX6OYKU>3,^8DW4@V+\_2A>9;gf:)
\A\<eL<&[K2;>S]UY,.JY[09F[bQS2@#BCPW?D<=#YTBVOf\DR/GPZaWTO8cQ@+c
#_aO<BL>[;@+Pg;/PWM+Q-XU#-gE<DX1GA4AgT[Y7G/:5SSK21c@dgFSD8=<5b8P
DF-]=S[-&S0g5[&47@0I_,Ybb3.1HZ;6:)UK2d4@^W+FSC5e#ggc\a#NVK?=SS;L
Ld=U,:L8Ab9D,T&GQ@cG3?bdAbPM<F2c;UO-FK224d8_:7X,7b#g<.PZ.K6+8+MB
K?Vbd5agG1XXP01#D@f]R/;LD13+2-O6&_\e<;_MGadDL1>g/)A(PeHdE231K3e0
&Z()IaR?bB6[VC\Y#Mf8]OagR(5W3)A[/ZUUC@1QWM20We\f.T-OeR7VQOWE2TSV
EA0(E,J9F_@P@cff7NY1>36.VQ&K<(GT?WZ.OWSBG5-V;dZg1@#>\X(D(2M9<15>
[\9Cg,X/cVf8\J;^_[-_?b4X<#,d&@R(0.JBFS0[V?_a3\^g3@Z[]fL]>G2R6YNV
F4/I0W,f[KFe<XS(c4G.CO/#_P4T]6+MS;U7W)];B(+=8K+)cfDe(c9U^^d,Z7<5
<[AF#</5OXNb3UJV.JG@/gHTVZe&K_CHB:1T.KM5<86)afAOMccI[1J4(MdSVXTC
2U)HGQbcd6A?a79Q@H>H?#@TOa\EKTG#0VfTE035Fb-;S-aQ-UaQJ@434XS#MP,T
T4H+NfC6A])Qc85aCU01=(1AXJ;dYQ:eGU7UMTDH,I][QXg;.8YEUKH4fgJW4XA.
EMeT_fMJ[d5K+QfM3:H37KAP_+f;aW29.&4+Pc.+;HD^?aY5:S]bX5?7b-b9=0ge
.U\WAY3bG1QN&@V&KU08aaS;KAe5\6^JR4:@+\_]H,V>5g[.R-BI1.<>,Ug2ffVK
E-A/+:SLXWM3=ZPSE#HEU^X7F-P>Q]J0U#UK?#O44U:O]GcQ/:Zgf1Q:S5QF&KG+
)<N(0;UVg7-fD>?eM<\Jd))>e#E&R[)@N?g>3&[Hb\b0fJ#U(<8)bT_CY/(]9&<?
LQ-<KWE.g8+Uc@FA&W7[EN7Ge4]cDQ;QJWQ30D:UX\QLNRgX1CD>HJbTNQP/QgHY
:XB0+?F)VKbE]ISHF2H)#E;=0I<c^dG6LER9gG]_>66HPTO2BN:UcDgf[2)Lg)C(
QN61T7>UB&:#G4^K#C0)JRCgU0P@@W]A=dW+&:49YU78GTe#G^aAT&R=4QZAT#9#
@e,]QZ1C7XQ<=#B\WSWIK6T^D._cCR4>GM(8U;7[@8/326_H;+5e6ASd3P:UKKZ]
eA0^PMK(MgA9b\2=PMcR<H:(RTG_/31+B5G7ZfT_-LNP-WXH-0[#>.]4L#ZRU30Q
W>fWWJ_=@+VW\7\Q5_O8Kf5H7N?8#;HdCL&,W#@BPO1^J&-;c)2c[CIaWXZ.6T5_
M(CT6b(V_XQ?/XGIO[R_6><fO_S=:>(YA4==#:K,J_G^9H1H?=3GN]Qf[6U8NX@V
->g65RF=6I<E[3[c.C.e_[>?)BV:\WPceR2U6K@QL2aa:8T/G>IRS;<O[9RD^<8I
_AeE:8U6f?SPAA_]D1<H&ZXA&=^\6WZC#gC>#g<P;NO)\J>Pa+YVAI\C0=Q^)75[
-Qc=4M08aR@5QUCA@GDfeO2J[+?ea^7b_C6X^3G^6N42@?C1D./:VH2#26S@M4]g
_,]eAe/aH]UK-2gO[DEaA&\TY-gLEC^8aS5+9a3MQQ.d)&I;]?QeUDQ5dP8&aL^C
;Mb/S0./S<&gMfY;UE81A0[7K]E9@e]b)aGISg9NYO6XeI8J<\1^OGZE51KNS>LX
7+<JYM_OBD?1fge23=e[12Y]HCY5Tb[@)3GF>2bA0K;fDUL0g6I80)Ib\=N8^6;a
TJ;D?Q(@>;f15K(TbdS-Q\f(,SdbWJYfeGT#(^7;BS&_2L=/BHf#K27?[@B5d_QC
I>/N-fM>3K:^V^R/c/_2LAN@C[NI8F7O<b#=-@Y78A#N]YM-2H4\L;)<eM<7Bb4Y
eM97:LFE@?,QKQ242EN4;bMI5HO_:cT4?^a-)I>BH/&>^;:7IFS(&Y4POTREgS1a
L(&#0TT<Z#S[G<1LRf-+>[a\[),X]T9O[DeX6@)PB;U=5Ug(;7&UG_=a34+1-01A
_XQ,&H@@gCMW\PcKEa<-XM\2ZI<D@44<9GFg3PK1Y^Pf(GJH];.a>=ZV@JP+/)DU
&Y3aLN6PN.=d@I4gaBZDI:^dUSaXT3P_LZJ/../e9N+W.-EV\QNE.+D\KI7NOP(I
&>JWe_XV=CTMO^+9]@fKfFYb4IcB=VA#JL[:<f,QgBPa(H.31Y41#OLbW77eY3_7
Ae6aDV#TN@=^>b(MQdWH[5K<Q8=E]3/bEGLNNf_(CJ<<SIP0:abXJT\0&\T@_)<:
5P)0MKP9EI90\KS_8@U.0/Df,&MS3:NJD)O<LM.]A+320R0>2fPBH^KM7W)?3f?Y
4?99d?CUFKJRUY=:Q^UbT]A@5RW.OI[DW7[c+dcH=U&EI<IB-:TIgI=LK#bIHQ96
/8FHJG52WID69W)SfA@0NY@:EKc1bHMBUY3\:2/GN8g2(MT7f@YUCB7B138eZ-P8
&^]9A+b9KXN83_DX<5.QRaNIW+^:)DBO@//0PS=d-U8EVIM8X;>=3:00]Pa5d9+M
e3I;PMSb[E[gf]c:eb(T6;9IKSJg6==ZV+I#AD3HT]4BgW#)ebH8)(X]3STaMG&(
C-4=)gX468.MBT#.a0#=)NBYJU,F8UDO[NP@N-A7c9SGHV=Rd-3>H(Zd)Z3a,g&d
T.^+fF4ab)&K7I2<M[=#,#,DUZF6]02,<8Odd&(+0L:D]OcM#>SGDAI2B?PC>J:V
BX9f?Ma^4aCIR27+:.W;K(QV&[JCb_QX:=Q4-#F&-ZEJ0Z/IBNg/5f,H13V&MgDV
dbG=4PVX;930)T^AAH<OGYB_Y3HYL_&A/&R5a#fJ22e;:<YCLX:V1[S)CAEd?(NT
,#>J8QdN57&eAXTG6OPSQ7G<RMIOKJ+T@X[RHJK8c#)fDLXYN4/DA42KQeE;CK9_
R^>9.I&Y(g@Ma58RbM67eVEY)0=Z]dWWK+98Z,]?KR1I4K@?gcZ3CUJ:5e,+&E>B
O/@,fNURaS=)(5=UZRfb-][I_Q[)YL>:EK(O_Ka@<=Y@K[O?2?92SBG[(9E[Ic)E
O1LRD8a^CS)G=.2I\2HVeGgeA#-C=1-[f<=d>MT\Fd(Q,@.DgH=/),04TOD,.<YB
O3Ke?:N>)cf\+9Ub=&S[>a(\KdT3Y7T7M:KL(d7&=]\-WE]OKD>4O\<0Cg?Te_\5
.5P#Ze+J0L6@R\b.U[\P8A/B#WA=ZB,[g+3((U4IPVD]CJ,\6PYOS@Z\4;Z8V?e)
94E>0.V?dNZR2VZN3X_I^NR[9?O^edRcR+UEf3&Q]@-gad2MfT0EV,FfW=FeP9c8
4:T=FZN_e8Z6FbTR3]4)YR++S+fP5<GTDNK^[AI#+->6K9#BJ+E^gFJ1\,,?;MA-
\.7.;d9[(.J&=2F_L_O@dU#eZ=5GWKMb&e7,[EG#X,V7SdeYB^MRgT1Y<IdHfK\(
[#/TdAP.JWF.A./JGNM34>^KBIQ]CEdW.Pf=:d(3@.#RdIQY[)d;]T?d#f4g_44M
2C,G=&VUR6^9U]?/(P.(BO^<bI?>8aIM>R0Q&U>Y=K&#(^1T3a@g_[^gc/@_JdY4
egQ>_e(2OT\1W,]#f-VTMFN_)/9+,Nf1R)LJbX>8IBXPa/ZE5USX053FI=BQ3gL,
DMVGE0&/58bM6J1N0Q<@a&IJ]?+.L+g(T\\c+U9)XPR3A2646d7_/+Bf5^d2H4-J
Q@-))B#V3dN8:&S6e#Z6/E#09VW@@MZIb4>28UY\e@GU+_Le2LM,<;>GOL_9YK2K
DW4CcL.QeZLF1,\+.(EK9AFWC9ebJ0X4ScWN9G6>=f1,FI(C\?](1C]3da^a<:E[
30WL[Ma^I&(-=?NS;&A_/eMDfYUWBM)O/7aC6U&=3#3P)a?S65IJA3@L@/@Z6Wd)
BUHO&0M[aZD)CWWAb<cVeN2ZEUDB\+C=)TOS\F=7@GG+V:0G@e#,.c7K=5E3IU]_
c#D1J+bKM^J5\EbO\:RL6.2[4BD0WK-f4g@](f4^W0dM7g10gS1@[V_DAN^6EC5G
KCfWa=IFHYg.;,@aba)f\8.=bTPCFfA/I:/_)Y)>DBR5@A(f;&>^YGg#@Y=I@AJ\
X.e1K,\O:]]\(.CN/&c73(Z28#9XQ;LFcUC3K-<aOd_gDX<L?Nb:BC_YVH,BEQ+G
+S;=PYKf9OO?c]3bZ=G=_O0QgIb2U4ff+0^0N;18?4#S=bVS@4a)[@2eQ&(E?a(]
8=50WfE2^ZFAYHM2+(EP.PE7Ee1C&H)^F68H1LI:Wf37eK=DBZP50+QZ7WB)SOK,
L&[P@Y.09J#3d>E&JZ5@.2[b3(B,Te;7b(3CF>MYB.Wa.X#KT>W#LH\#[0TE22M.
K\/UM3_^IHfaF9HSZ5,@;+@7PN^:\)\0L+_Xf0CcIG/?),@(9O.f.:5IIF](g55@
TR_9KVe3L^9f^S-2G6UJTU:KQFd&YA]LEQT1@T^M:/;2BdUY6H>E83F_.4/PY[K^
@JAJ>S(Z0@]3P,@G9E[X]&CT:@TeHe1DTKfg9V)N4)PL:D/g(F2_U@3Z&2CAaBW.
R=Qg+XNMH;B7S4F?8fU0^gc7I.a,(P^C/\?1)&;;Q]#AVTAA,(6NQ4S(8HJ6YX1B
JV+WW[+EQVT/N,e-+[bW7#DBQ\TZ?]V09J)UHG+5TXM1R2fI4R>>,0&a?-YIP/<?
YQ:g?<6</&XVMKG,]UZ(SU=FO;61W<2E718VKCXNS,IQ1_]<IX#2-1BP9:J\V,bd
.1a-8Y(gHc2YXM+NSF20_AMQJGIJDK6b_I+G+^F=Q&34BgQ+\,^7.KXWLU[>0#W3
4dAHW^5<S.8JCf]2JW=4W@MQ\0LZQa==4UcH&FG8OgRHJ)8+D#&gJc=M[cD.SdM@
QRG3DB&V.4;;2&3_=\P5+GOUGMW+9RdZ7PZ4@;&ETO.I/M9))b3=_d.U>>5@)(]Y
H61,G17J1QFQQGae93[RcUR6FUF:8(=e[V(fR?#E[6#GRW^C@NQG_<W[2gG(#5b6
U@cPK]YZG5\bOgJ8_:B6RGaI#C<F>G79>3-41Bb1,FC1#?G.[>5b3TX=>M(QgD8U
a&PR:@,2;6TROLU7[gB3d^X0SR=_f6eFB3fd>YNc65:eBdZK.W364XdK1ZQ-,:/Y
(?V]Q4PEYG<:I-UaIXN54JCXc/Z@ZKX-gH,85KBCdIY[L,NI;3b.a7V7)@_-6JZC
E<G9KR6I-PXX1N0RM8XXTHCX3$
`endprotected


ps p(bif.TI,bif.FO);

initial begin
//    repeat(10_000_000) @(posedge(clk));
    $dumpfile("perm.vcd");
    $dumpvars(9,top);
    repeat(100000) @(posedge(clk));
    #5;
    $dumpoff;

end

endmodule : top
